//--------------------------------------------------------------------------------
//  %file% - Time-stamp: <Sat Dec 22 12:29:55 JST 2018>
//
//   Copyright (c) %year%  %id% (%name%)  <%mail%>
//
//  $Id: %file% %date% %id% $
// Create Date: %date%
// Design Name:
// Module Name: %file%
// Project Name: 
// Target Devices:
// Tool versions:
// Description: 
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//--------------------------------------------------------------------------------

module modulename #(parameter WIDTH= 8)
   (
    input wire 			   clk,
    input wire 			   rst,
	output wire 		   out1,
	output reg [WIDTH-1:0] out2
    );
   
endmodule // modulename
